module can_rx
#(
	parameter smth = 0
)(
	input rst_i,
	input clk_can_i
);
reg as;


endmodule 